/** 
 * @info    Testbench for the SIMON top module
 * 
 * @author Anastasios Psarras (a.psarras4225@gmail.com)
 *
 * @license MIT license, check license.md
 * 
 * @brief -- To run the testbench you need a simulator that supports SystemVerilog & DPI-C:
 *           1. Compile files contained in <./flist>
 *           2. Simulate & run
 *              Your output should be flooded with *** INFO *** and *** SUCCESS *** messages,
 *              ending with: [chck] *** INFO *** Checked all transactions: 100/100 succeeded.
 *              If you get less than 100% verified transactions, something has gone wrong.
 *              Make sure your simulator breaks on Error, so that you don't miss possible errors.
 *
 *        -- To customize the RTL:
 *           To generate and run any Simon 2n/mn configuration, set parameters WW and NKW  accordingly,
 *           where n=WW (word size), and m=NKW (key size). Default values are WW=32, NKW=3, which generates Simon 64/96.
 *           Note that the verification environment only supports Simon 64/96, 64/128, 128/128, 128/192, 128/256,
 *           since NSA provides reference C code only for those configurations. RTL supports all possible configurations.
 *
 *        -- To customize the TB:
 *           You can change the number of random transactions generated by setting ITEMS_TO_GENERATE parameter in tb_top.
 *           Each transaction is randomly selected to be an encryption or decryption process, in which case, a random Default
 *           value is 100, i.e. 100 random plaintext-key or ciphertext-key pairs are generated.
 *
 */
 
`timescale 1ps/1ps

// `default_nettype none
module tb_top
#(
)
(
);

// -- Imports ------------------------------------------------------------------------------------- //
import tb_crypto_item_pkg::crypto_item;
import simon_const_pkg::*;
import "DPI-C" function void dpi_c_run_simon(input int crypto_mode, byte txt_i[], byte key_i[], output byte txt_o[]);

/*       Manual ENC | DEC | Auto
 32-3:          OK  | OK  |  OK
 32-4:          OK  | OK  |  OK
 64-2:          OK  | OK  |  OK
 64-3:          OK  | OK  |  OK
 64-4:          OK  | OK  |  OK
*/

// -- RTL Config ---------------------------------------------------------------------------------- //
localparam int   WW                 = 64;
localparam int   NKW                = 3;
localparam logic DATA_RST           = 1'b0;
// -- TB Config ----------------------------------------------------------------------------------- //
localparam int   ITEMS_TO_GENERATE  = 100;

// -- clk/rst ------------------------------------------------------------------------------------- //
localparam CLK_PERIOD = 200;
logic clk, arst_n;
    
initial begin clkrst:
    clk = 0;
    arst_n = 1;
    #(CLK_PERIOD/2) arst_n = 0;
    #(2*CLK_PERIOD+CLK_PERIOD/2) arst_n = 1;
end
always #(CLK_PERIOD/2) clk = ~clk;

// -- DUT ----------------------------------------------------------------------------------------- //
logic                    active_o;
logic                    simon_inp_valid;
logic                    simon_inp_ready;
logic                    simon_inp_mode;
logic[2-1:0][WW-1:0]     simon_inp_pt;
logic[NKW-1:0][WW-1:0]   simon_inp_key;
logic                    simon_out_valid;
logic                    simon_out_ready;
logic                    simon_out_mode;
logic[2-1:0][WW-1:0]     simon_out_ct;

simon_top
#(
    .WW             (WW),
    .NKW            (NKW),
    .DATA_RST       (DATA_RST)
)
i_core
(
    .clk            (clk),
    .arst_n         (arst_n),
    
    .active_o       (active_o),
    
    .valid_i        (simon_inp_valid),
    .ready_o        (simon_inp_ready),
    .mode_i         (simon_inp_mode),
    .pt_i           (simon_inp_pt),
    .key_i          (simon_inp_key),
    
    .valid_o        (simon_out_valid),
    .ready_i        (simon_out_ready),
    .mode_o         (simon_out_mode),
    .ct_o           (simon_out_ct)
);

// -- Interface with SIMON ------------------------------------------------------------------------ //
task automatic write_to_input(input logic mode, logic[2-1:0][WW-1:0] pt, logic[NKW-1:0][WW-1:0] key);
    simon_inp_valid   <= 1;
    simon_inp_mode    <= mode;
    simon_inp_pt      <= pt;
    simon_inp_key     <= key;
    
    do begin
        @(posedge clk);
    end while (!simon_inp_ready);
    
    simon_inp_valid   <= 0;
    simon_inp_mode    <= 'x;
    simon_inp_pt      <= 'x;
    simon_inp_key     <= 'x;
endtask

// blocking read from output
task automatic read_from_output_b(ref logic[2-1:0][WW-1:0] ct, logic mode);
    simon_out_ready <= 1;
    
    do begin
        @(posedge clk);
    end while (!simon_out_valid);
    ct  = simon_out_ct;
    mode = simon_out_mode;
    simon_out_ready <= 0;
endtask

// -- Mailboxes ----------------------------------------------------------------------------------- //
mailbox #(crypto_item #(.WW(WW), .NKW(NKW) )) mb_source_2_driver;
mailbox #(crypto_item #(.WW(WW), .NKW(NKW) )) mb_driver_2_checker;
mailbox #(crypto_item #(.WW(WW), .NKW(NKW) )) mb_sink_2_checker;

// -- TB ------------------------------------------------------------------------------------------ //
initial begin
    mb_source_2_driver = new();
    mb_driver_2_checker = new();
    mb_sink_2_checker = new();
    
    @(negedge arst_n);
    @(posedge arst_n);
    $display("%0t: [mngr] *** INFO *** Reset phase ended.", $time);
    
    fork
        do_source();
        do_driver();
        do_sink();
        do_checker();
    join_none
    $display("%0t: [mngr] *** INFO *** Started everything.", $time);
end

// -- Source -------------------------------------------------------------------------------------- //
task automatic do_source();
    for (int i=0; i<ITEMS_TO_GENERATE; i++) begin
        crypto_item #(.WW(WW), .NKW(NKW) ) the_item;
        
        @(posedge clk);
        // Produce a random item
        the_item                = new();
        assert (the_item.randomize()) else $error("Failed to randomize item");
        
        // the_item.crypto_mode    = MODE_DEC;
        // the_item.txt            = '{8'h_72, 8'h_69, 8'h_62, 8'h_65, 8'h_20, 8'h_77, 8'h_68, 8'h_65, 8'h_6e, 8'h_20, 8'h_74, 8'h_68, 8'h_65, 8'h_72, 8'h_65, 8'h_20};
        // the_item.key            = '{8'h_00, 8'h_01, 8'h_02, 8'h_03, 8'h_04, 8'h_05, 8'h_06, 8'h_07, 8'h_08, 8'h_09, 8'h_0a, 8'h_0b, 8'h_0c, 8'h_0d, 8'h_0e, 8'h_0f, 8'h_10, 8'h_11, 8'h_12, 8'h_13, 8'h_14, 8'h_15, 8'h_16, 8'h_17};
        // the_item.txt            = '{8'h_5b, 8'h_b8, 8'h_97, 8'h_25, 8'h_6e, 8'h_8d, 8'h_9c, 8'h_6c, 8'h_4f, 8'h_0d, 8'h_dc, 8'h_fc, 8'h_ef, 8'h_61, 8'h_ac, 8'h_c4};

        the_item.gen_time = $time();
        // Push to [Source]-->[Driver] mailbox
        assert (mb_source_2_driver.try_put(the_item)) else $error("[Source] could not put int mb_source_2_driver");
        $display("%0t: [srce] *** INFO *** produced item:\n      %s", $time, the_item.to_str(the_item.crypto_mode == MODE_ENC));
    end
    $display("%0t: [srce] *** INFO *** ended production of %0d items", $time, ITEMS_TO_GENERATE);
endtask
/*
64/96
    the_item.txt            = '{8'h_63, 8'h_6c, 8'h_69, 8'h_6e, 8'h_67, 8'h_20, 8'h_72, 8'h_6f};
    the_item.key            = '{8'h_00, 8'h_01, 8'h_02, 8'h_03, 8'h_08, 8'h_09, 8'h_0a, 8'h_0b, 8'h_10, 8'h_11, 8'h_12, 8'h_13};
    the_item.txt            = '{8'h_c8, 8'h_8f, 8'h_1a, 8'h_11, 8'h_7f, 8'h_e2, 88'h_a2, 8'h_5c};
64/128
    the_item.txt            = '{8'h_75, 8'h_6e, 8'h_64, 8'h_20, 8'h_6c, 8'h_69, 8'h_6b, 8'h_65};
    the_item.key            = '{8'h_00, 8'h_01, 8'h_02, 8'h_03, 8'h_08, 8'h_09, 8'h_0a, 8'h_0b, 8'h_10, 8'h_11, 8'h_12, 8'h_13, 8'h_18, 8'h_19, 8'h_1a, 8'h_1b};
    the_item.txt            = '{8'h_7a, 8'h_a0, 8'h_df, 8'h_b9, 8'h_20, 8'h_fc, 8'h_c8, 8'h_44};
128/128
    the_item.txt            = '{8'h_20, 8'h_74, 8'h_72, 8'h_61, 8'h_76, 8'h_65, 8'h_6c, 8'h_6c, 8'h_65, 8'h_72, 8'h_73, 8'h_20, 8'h_64, 8'h_65, 8'h_73, 8'h_63};
    the_item.key            = '{8'h_00, 8'h_01, 8'h_02, 8'h_03, 8'h_04, 8'h_05, 8'h_06, 8'h_07, 8'h_08, 8'h_09, 8'h_0a, 8'h_0b, 8'h_0c, 8'h_0d, 8'h_0e, 8'h_0f};
    the_item.txt            = '{8'h_bc, 8'h_0b, 8'h_4e, 8'h_f8, 8'h_2a, 8'h_83, 8'h_aa, 8'h_65, 8'h_3f, 8'h_fe, 8'h_54, 8'h_1e, 8'h_1e, 8'h_1b, 8'h_68, 8'h_49};
128/192
    the_item.txt            = '{8'h_72, 8'h_69, 8'h_62, 8'h_65, 8'h_20, 8'h_77, 8'h_68, 8'h_65, 8'h_6e, 8'h_20, 8'h_74, 8'h_68, 8'h_65, 8'h_72, 8'h_65, 8'h_20};
    the_item.key            = '{8'h_00, 8'h_01, 8'h_02, 8'h_03, 8'h_04, 8'h_05, 8'h_06, 8'h_07, 8'h_08, 8'h_09, 8'h_0a, 8'h_0b, 8'h_0c, 8'h_0d, 8'h_0e, 8'h_0f, 8'h_10, 8'h_11, 8'h_12, 8'h_13, 8'h_14, 8'h_15, 8'h_16, 8'h_17};
    the_item.txt            = '{8'h_5b, 8'h_b8, 8'h_97, 8'h_25, 8'h_6e, 8'h_8d, 8'h_9c, 8'h_6c, 8'h_4f, 8'h_0d, 8'h_dc, 8'h_fc, 8'h_ef, 8'h_61, 8'h_ac, 8'h_c4};
128/256
    the_item.txt            = '{8'h_69, 8'h_73, 8'h_20, 8'h_61, 8'h_20, 8'h_73, 8'h_69, 8'h_6d, 8'h_6f, 8'h_6f, 8'h_6d, 8'h_20, 8'h_69, 8'h_6e, 8'h_20, 8'h_74};
    the_item.key            = '{8'h_00, 8'h_01, 8'h_02, 8'h_03, 8'h_04, 8'h_05, 8'h_06, 8'h_07, 8'h_08, 8'h_09, 8'h_0a, 8'h_0b, 8'h_0c, 8'h_0d, 8'h_0e, 8'h_0f, 8'h_10, 8'h_11, 8'h_12, 8'h_13, 8'h_14, 8'h_15, 8'h_16, 8'h_17, 8'h_18, 8'h_19, 8'h_1a, 8'h_1b, 8'h_1c, 8'h_1d, 8'h_1e, 8'h_1f};
    the_item.txt            = '{8'h_68, 8'h_b8, 8'h_e7, 8'h_ef, 8'h_87, 8'h_2a, 8'h_f7, 8'h_3b, 8'h_a0, 8'h_a3, 8'h_c8, 8'h_af, 8'h_79, 8'h_55, 8'h_2b, 8'h_8d};
*/

// -- Driver -------------------------------------------------------------------------------------- //
task automatic do_driver();
    simon_inp_valid <= 0;
    simon_inp_mode  <= 'x;
    simon_inp_pt    <= 'x;
    simon_inp_key   <= 'x;
    // start driver loop
    forever begin
        crypto_item #(.WW(WW), .NKW(NKW) ) the_item;
        logic[2-1:0][WW-1:0]    the_txt;
        logic[NKW-1:0][WW-1:0]  the_key;
        
        @(posedge clk);
        // -- Mailbox Read -- //
        mb_source_2_driver.get(the_item);
        $display("%0t: [drvr] *** INFO *** got item from mb:\n      %s", $time, the_item.to_str(the_item.crypto_mode == MODE_ENC));
        
        the_txt = the_item.get_word_packed_txt();
        the_key = the_item.get_word_packed_key();
        $display("%0t: [drvr] *** INFO *** driving pt: %h %h | key: %h", $time, the_txt[1], the_txt[0], the_key);
        
        if (the_item.crypto_mode == MODE_DEC) begin
            the_txt = {the_txt[0], the_txt[1]}; // word reverse!
        end
        write_to_input(.mode(the_item.crypto_mode), .pt(the_txt), .key(the_key));
        assert (mb_driver_2_checker.try_put(the_item)) else $error("[drvr] *** ERROR *** could not put int mb_driver_2_checker");
    end
endtask

// -- Sink ---------------------------------------------------------------------------------------- //
task automatic do_sink();
    simon_out_ready <= 0;
    
    // start sink loop
    forever begin
        logic[2-1:0][WW-1:0]    the_txt;
        logic                   the_mode;
        crypto_item #(.WW(WW), .NKW(NKW) ) the_item;
        
        @(posedge clk);
        read_from_output_b(the_txt, the_mode);
        the_item                = new();
        the_item.key            = '{NKW*WW/8{8'b0}};
        the_item.crypto_mode    = the_mode;
        if (the_mode == MODE_DEC) begin
            the_txt = {the_txt[0], the_txt[1]};
        end
        the_item.set_txt_from_packed_words(the_txt);
        
        $display("%0t: [sink] *** INFO *** got item from simon:\n      %s", $time, the_item.to_str(the_item.crypto_mode == MODE_DEC));
        assert (mb_sink_2_checker.try_put(the_item)) else $error("[sink] *** ERROR *** could not put int mb_sink_2_checker");
    end
endtask

// -- Checker ------------------------------------------------------------------------------------- //
task automatic do_checker();
    automatic int total_count = 0;
    automatic int success_count = 0;
    
    while (total_count < ITEMS_TO_GENERATE) begin
        crypto_item #(.WW(WW), .NKW(NKW) ) item_in;
        crypto_item #(.WW(WW), .NKW(NKW) ) item_out;
        crypto_item #(.WW(WW), .NKW(NKW) ) item_gold;
        
        // Read from mailboxes for new items -- blocking reads
        mb_driver_2_checker.get(item_in);
        mb_sink_2_checker.get(item_out);
        
        $display("%0t: [chck] *** INFO *** got source item: %s", $time, item_in.to_str(item_in.crypto_mode == MODE_ENC));
        $display("%0t: [chck] *** INFO *** got sink item:   %s", $time, item_out.to_str(item_out.crypto_mode == MODE_DEC));
        
        if (item_in.crypto_mode == item_out.crypto_mode) begin
            byte golden_txt[2*WW/8];
            $display("%0t: [chck] *** INFO *** Calling DPI-C golden routine for %scryption...", $time, item_in.crypto_mode == MODE_ENC ? "en" : "de");
            dpi_c_run_simon(.crypto_mode(int'(item_in.crypto_mode)), .txt_i(item_in.txt), .key_i(item_in.key), .txt_o(golden_txt));
            item_gold = new();
            item_gold.txt = golden_txt;
            if (golden_txt == item_out.txt) begin
                success_count++;
                $display("%0t: [chck] *** SUCCESS *** Generated (%s) matches Golden (%s)", $time, item_out.txt_to_str(), item_gold.txt_to_str());
            end else begin
                $error("%0t: [chck] *** FAILURE *** Generated (%s) does NOT match Golden (%s)", $time, item_out.txt_to_str(), item_gold.txt_to_str());
            end
        end else begin
            $error("%0t: [chck] *** FAILURE *** source/sink items' << MODE >> DO NOT match! ", $time);
        end
        
        total_count++;
    end
    
    $display("\n");
    $display("%0t: [chck] *** INFO *** Checked all transactions: %0d/%0d succeeded.", $time, success_count, total_count);
    $display("\n");
    $display("%0t: [chck] *** INFO *** Now ending", $time);
    $display("\n");
    $finish();
endtask


endmodule
// `default_nettype wire