/**
 * @info Package containing SIMON constants
 *
 * @author Anastasios Psarras (a.psarras4225@gmail.com)
 *
 * @license MIT license, check license.md
 *
 */

package simon_const_pkg;

localparam logic MODE_ENC = 1'b0;
localparam logic MODE_DEC = 1'b1;

endpackage